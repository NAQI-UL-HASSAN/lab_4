module RGBLAB_tb();
    logic a0, a1, b0, b1, R1, G1, B1;
    RGBLAB DUT(
        .a_0(a0),
        .a_1(a1),
        .b_0(b0),
        .b_1(b1),
        .R(R1),
        .G(G1),
        .B(B1)
    );
    initial
    begin
    a0 = 0; a1 = 0; b0 = 0; b1 = 0;
    #10;
    a0 = 0; a1 = 0; b0 = 0; b1 = 1;
    #10;
    a0 = 0; a1 = 0; b0 = 1; b1 = 0;
    #10;
    a0 = 0; a1 = 0; b0 = 1; b1 = 1;
    #10;
    a0 = 0; a1 = 1; b0 = 0; b1 = 0;
    #10;
    a0 = 0; a1 = 1; b0 = 0; b1 = 1;
    #10;
    a0 = 0; a1 = 1; b0 = 1; b1 = 0;
    #10;
    a0 = 0; a1 = 1; b0 = 1; b1 = 1;
    #10;
    a0 = 1; a1 = 0; b0 = 0; b1 = 0;
    #10;
    a0 = 1; a1 = 0; b0 = 0; b1 = 1;
    #10;
    a0 = 1; a1 = 0; b0 = 1; b1 = 0;
    #10;
    a0 = 1; a1 = 0; b0 = 1; b1 = 1;
    #10;
    a0 = 1; a1 = 1; b0 = 0; b1 = 0;
    #10;
    a0 = 1; a1 = 1; b0 = 0; b1 = 1;
    #10;
    a0 = 1; a1 = 1; b0 = 1; b1 = 0;
    #10;
    a0 = 1; a1 = 1; b0 = 1; b1 = 1;
    #10;
    $stop;   
    end
endmodule